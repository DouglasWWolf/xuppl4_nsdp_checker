
//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 27-Apr-2024  1.0.0  DWW  Initial creation
//================================================================================================
localparam RTL_TYPE      = 12266;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 27;
localparam VERSION_MONTH = 4;
localparam VERSION_YEAR  = 2024;

/*
================================================================================================
  Vers      Date      Who  Changes
 -----------------------------------------------------------------------------------------------
  1.0.0  27-Apr-2024  DWW  Initial creation
                                                   
  1.1.0  04-May-2024  DWW  Now checking RDMX target addresses in the packet headers
                                                      
  1.2.0  21-May-2024  DWW  Now ignoring sensor-chip frame-header cells when checking frame-data
                           for correctness.
                                                         
  1.3.0  22-May-2024  DWW  Made the logic that ignores sensor-chip frame-headers aware of 
                           "PACKETS_PER_GROUP".  This is because the number of packets with 
                           sensor-chip headers that each channel sees depends on the number of
                           packets per ping-pong group.
                                                           
  1.4.0  22-May-2024  DWW  Added logic to ignore sensor-chip frame-footers

  2.1.0  19-Jun-2025  DWW  Integration with new build/release system
                           Added check for sender's QSFP port
                           Added check for RDMX flags 
================================================================================================
*/

localparam RTL_TYPE      = 12266;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_MAJOR = 2;
localparam VERSION_MINOR = 1;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;


//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 27-Apr-2024  1.0.0  DWW  Initial creation
//
// 04-May-2024  1.1.0  DWW  Now checking RDMX target addresses in the packet headers
//
// 21-May-2024  1.2.0  DWW  Now ignoring senor-chip frame-header cells when checking frame-data
//                          for correctness.
//================================================================================================
localparam RTL_TYPE      = 12266;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 2;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 21;
localparam VERSION_MONTH = 5;
localparam VERSION_YEAR  = 2024;
